

module sqeuential {
	input  CLOCK_50,

	input [3:0] KEY,

	output [9:0] LEDR,

	input [9:0] SW

};

endmodule

module parallel_load(input btn, clk, input [4:0] in, output [4:0] out);

endmodule
